module top_bridge ();


endmodule

module mac1100 ();
Triple_Speed_Ethernet_MAC_Top mac1100 ();

//TODO()
endmodule

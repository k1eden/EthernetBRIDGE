module txfifo ();

//TODO()
endmodule

module mac1200 ();

//TODO()
endmodule

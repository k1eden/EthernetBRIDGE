module rxfifo ();

//TODO()
endmodule

module mac1100 ();

//TODO()
endmodule
